module adyacentes(input clk, input logic [7:0][7:0] matriz, input logic[1:0] celda);


endmodule
