module minesweeper(
);

endmodule